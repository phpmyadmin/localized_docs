PO4A-HEADER:mode=before;position=<head>
<!--

Denna fil skapas med hjälp av po4a, editera ej!

Du kan redigera po filer för att ändra översättningen.

Eller så kan du redigera dom via internet på
https://l10n.cihar.com/projects/pmadoc/.

-->
